module repo_template

pub fn hello() string {
	return 'Hello World'
}
